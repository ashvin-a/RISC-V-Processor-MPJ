/////////////////////////////////////////////////////////////
///////////////////////// HAZARD CONTROL UNIT////////////////////
/////////////////////////////////////////////////////////////

module hazard_control_unit();
endmodule